** Profile: "SCHEMATIC1-t"  [ c:\users\hp\documents\tencent files\740167442\filerecv\temperature_1pspice\temperature_1\t-pspicefiles\schematic1\t.sim ] 

** Creating circuit file "t.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
.INC "c:\users\hp\documents\tencent files\740167442\filerecv\temperature_1pspice\temperature_1\t-pspicefiles\schematic1\t\t_profile"
+ ".inc" 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 20m 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
