** Profile: "SCHEMATIC1-w3"  [ C:\Workspace\Cadence\01\w3-pspicefiles\schematic1\w3.sim ] 

** Creating circuit file "w3.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5ms 1u 1u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
